module New_module();

endmodule : New_module