package New_package;
// why do all bands now sound like pop shit?
// another pull test, how will deleting and recreating document look?
endpackage
