module New_module_sv();

endmodule : New_module_sv