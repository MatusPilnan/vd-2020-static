module New_module();
//changed
endmodule : New_module