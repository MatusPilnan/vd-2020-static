package New_package;
// why do all bands now sound like pop shit?
// tried to change that?
endpackage
