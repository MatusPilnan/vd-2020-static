package New_package;
// why do all bands now sound like pop shit?
// will it work from app?
// be a conflict
endpackage
