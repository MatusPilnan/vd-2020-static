package New_package;

endpackage