module New_module();
//changed
// now there should be an actual commit message
endmodule : New_module