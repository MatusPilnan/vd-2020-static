module aj_toto_by_som_skusil_sv();

endmodule : aj_toto_by_som_skusil_sv