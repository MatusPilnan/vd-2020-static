package New_package;
// why do all bands now sound like pop shit?
// now with op?
endpackage
